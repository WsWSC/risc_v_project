//////////////////////////////////////////////////
// risc v side project                          //
//                                              //
// create by WsWSC                              //
//////////////////////////////////////////////////

module regs(
    input wire clk,
    input wire rst,

    // from id
    input wire[4:0]     reg1_raddr_i,
    input wire[4:0]     reg2_raddr_i,

    // to id
    output reg[31:0]    reg1_rdata_o,
    output reg[31:0]    reg2_rdata_o,

    // from ex
    input wire[4:0]     reg_waddr_i,
    input wire[31:0]    reg_wdata_i,
    input               reg_wen
);

    reg[31:0] regs[0:31];
    integer i;              // initial for loop

    // id stage, read rs1 data
    always@(*) begin
        if(rst == 1'b0) 
            reg1_rdata_o <= 32'b0;
        else if (reg1_raddr_i == 5'b0)
            reg1_rdata_o <= 32'b0;
        else if (reg_wen && (reg_1_raddr_i == reg_waddr_i) )    // hazard detection
            reg1_rdata_o <= reg[reg1_raddr_i];
        else 
            reg1_rdata_o <= regs[reg1_raddr_i];
    end

    // id stage, read rs2 data
    always@(*) begin
        if(rst == 1'b0) 
            reg2_rdata_o <= 32'b0;
        else if (reg2_raddr_i == 5'b0)
            reg2_rdata_o <= 32'b0;
        else if (reg_wen && (reg_2_raddr_i == reg_waddr_i) )    // hazard detection
            reg2_rdata_o <= reg[reg2_raddr_i];
        else 
            reg2_rdata_o <= regs[reg2_raddr_i];
    end

    // ex stage, wirte reg 
    always@(posedge clk) begin
        if(rst == 1'b0) begin
            for (i = 1; i <= 31; i = i + 1) begin     // reg x0 is always 0, no need reset
                reg[i] <= 32'b0;
            end
        end else 
            reg[reg_waddr_i] <= reg_wdata_i;
    end

endmodule