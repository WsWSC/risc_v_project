module top(
    input wire clk,
    input wire rst_n,
    input wire [31:0] inst_i,

    output wire [31:0] inst_addr_o
);




endmodule